library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DeCoder is
    Port ( selector : in  STD_LOGIC_VECTOR (4 downto 0);
			  reg : out  STD_LOGIC_VECTOR (31 downto 0);
			  E:IN  STD_LOGIC );
		
end DeCoder;

architecture Behavioral of DeCoder is

begin
reg <= "00000000000000000000000000000000"	WHEN E = '0' ELSE
"00000000000000000000000000000001" WHEN selector = "00000" ELSE
"00000000000000000000000000000010" WHEN selector = "00001" ELSE
"00000000000000000000000000000100" WHEN selector = "00010" ELSE
"00000000000000000000000000001000" WHEN selector = "00011" ELSE
"00000000000000000000000000010000" WHEN selector = "00100" ELSE
"00000000000000000000000000100000" WHEN selector = "00101" ELSE
"00000000000000000000000001000000" WHEN selector = "00110" ELSE
"00000000000000000000000010000000" WHEN selector = "00111" ELSE
"00000000000000000000000100000000" WHEN selector = "01000" ELSE
"00000000000000000000001000000000" WHEN selector = "01001" ELSE
"00000000000000000000010000000000" WHEN selector = "01010" ELSE
"00000000000000000000100000000000" WHEN selector = "01011" ELSE
"00000000000000000001000000000000" WHEN selector = "01100" ELSE
"00000000000000000010000000000000" WHEN selector = "01101" ELSE
"00000000000000000100000000000000" WHEN selector = "01110" ELSE
"00000000000000001000000000000000" WHEN selector = "01111" ELSE
"00000000000000010000000000000000" WHEN selector = "10000" ELSE
"00000000000000100000000000000000" WHEN selector = "10001" ELSE
"00000000000001000000000000000000" WHEN selector = "10010" ELSE
"00000000000010000000000000000000" WHEN selector = "10011" ELSE
"00000000000100000000000000000000" WHEN selector = "10100" ELSE
"00000000001000000000000000000000" WHEN selector = "10101" ELSE
"00000000010000000000000000000000" WHEN selector = "10110" ELSE
"00000000100000000000000000000000" WHEN selector = "10111" ELSE
"00000001000000000000000000000000" WHEN selector = "11000" ELSE
"00000010000000000000000000000000" WHEN selector = "11001" ELSE
"00000100000000000000000000000000" WHEN selector = "11010" ELSE
"00001000000000000000000000000000" WHEN selector = "11011" ELSE
"00010000000000000000000000000000" WHEN selector = "11100" ELSE
"00100000000000000000000000000000" WHEN selector = "11101" ELSE
"01000000000000000000000000000000" WHEN selector = "11110" ELSE
"10000000000000000000000000000000" WHEN selector = "11111" ;

end Behavioral;